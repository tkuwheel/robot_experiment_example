library verilog;
use verilog.vl_types.all;
entity halfadd_vlg_vec_tst is
end halfadd_vlg_vec_tst;
